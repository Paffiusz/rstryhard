
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity emitter is
end emitter;

architecture Behavioral of emitter is

begin


end Behavioral;

